�� sr java.util.ArrayListx����a� I sizexp   w   sr com.sut.parpar.Player��I�;�.� Z 
cutterFLAGZ 	isSpeedupZ 	isgodMODEI playerIDI powerupSTARTZ 	splitFLAGJ 	splitTimeI tickD velXD velYL biggestCirlet )Lcom/sut/parpar/gameobjects/MovingCircle;L circlest Ljava/util/ArrayList;L imaget Ljava/awt/image/BufferedImage;L namet Ljava/lang/String;L playerColort Ljava/awt/Color;L powerUpt $Lcom/sut/parpar/gameobjects/PowerUp;L spawnert Lcom/sut/parpar/Spawner;xp                �  t                sr 'com.sut.parpar.gameobjects.MovingCircle%��3�p Z isEatenZ isGodZ isSpeedI playerIDL spawnerq ~ 	xr !com.sut.parpar.gameobjects.Circlel�i�R��  xr %com.sut.parpar.gameobjects.GameObjectUP,\*I 	D radiusD surfaceD velXD velYD widthD xD yL colorq ~ L typet 'Lcom/sut/parpar/gameobjects/ObjectType;xp@,"Vl�@�Y���#Y�\8��P�@X�b��@<"Vl�@�s�b$�n@�%^���sr java.awt.Color���3u F falphaI valueL cst Ljava/awt/color/ColorSpace;[ 	frgbvaluet [F[ fvalueq ~ xp    ��  ppp~r %com.sut.parpar.gameobjects.ObjectType          xr java.lang.Enum          xpt PLAYER      sr com.sut.parpar.Spawner�&�� �� I heightI maxNumofFoodI widthL foodsq ~ L powerUpq ~ L sawt  Lcom/sut/parpar/gameobjects/Saw;xp  \     �sq ~     w   sr com.sut.parpar.gameobjects.Food�X.	�Q Z isEatenxq ~ ?�^E!ZM@&������                @^E!ZM@\�&�H9�@l_��
g"sq ~     �ߜ�ppp~q ~ t ORDINARY_FOOD sq ~ @$"�>�|N@s�ν��                @4"�>�|N@�тmM4�@gR��8�sq ~     �fZpppq ~  sq ~ @*G�Ϻ�@��N�u                @:G�Ϻ�@���7�@��Hz�psq ~     ��pppq ~  sq ~ @&�k�M��@y�T��P                @6�k�M��@������@|5�:��sq ~     ��ֿpppq ~  sq ~ @"���@p��bi�                @2���@�-��G#�@{�a�	�sq ~     �n�,pppq ~  sq ~ @��"	�@i;x�F                @/��"	�@����0�@b:7���8sq ~     ���pppq ~  sq ~ @"hq�g@p��P�,                @2hq�g@n-9���@v%�*F+sq ~     �K��pppq ~  sq ~ @#.P���_@rC��?�                @3.P���_@n
IH�!�@v�@7g�sq ~     ��vpppq ~  sq ~ @,%~Wo�K@�q�V �                @<%~Wo�K@�P�Yw�@{҆�Q�sq ~     ��V^pppq ~  sq ~ @���9@]u���5                @(���9@���5 �@u@�H���sq ~     ����pppq ~  sq ~ ?�4��2.t@$�p!�V_                @4��2.t@z鷏�#@w�ؚC�2sq ~     �il�pppq ~  sq ~ @({�ο�7@}lx�ݚ�                @8{�ο�7@��&�P%�@r�˳���sq ~     �%pppq ~  sq ~ @*>�w��@���@�                @:>�w��@r���~�@Z��nsq ~     �2�pppq ~  sq ~ ?�n�saڲ?�N��q                ?�n�saڲ@���+�@\��U�xsq ~     �?؟pppq ~  sq ~ @(K�>f�@|�U��                @8K�>f�@z"ik�@��ߴ��sq ~     �^� pppq ~  sq ~ @'+����@z[T}Oٝ                @7+����@�{��@xM.���sq ~     � �pppq ~  sq ~ @��QF�@c	��Fp^                @+��QF�@�i��(�@�I�4/(sq ~     �mK�pppq ~  sq ~ @.L��@<�9�Pt                @.L��@�}je�1@�@L�u�sq ~     �H�pppq ~  sq ~ @"��&@qw��`�                @2��&@�Z���%�@��=�g�sq ~     �C�pppq ~  sq ~ @����7@iӻ��=                @/����7@���P�#�@����Sf�sq ~     �u��pppq ~  sq ~ @#�Q�?��@s\�ׁN2                @3�Q�?��@��KyN��@v�#�sq ~     �:܂pppq ~  xsr "com.sut.parpar.gameobjects.PowerUp�5����F  xq ~                                 @4      @�[�Y]�@�9�|�0sq ~     ��&.ppp~q ~ t GOD_MODE sr com.sut.parpar.gameobjects.SawB�z�b I scalexq ~                                 @T      @�]�qj@r{�ۍ��sq ~     �ΐbppp~q ~ t SAW    sq ~     w   sq ~ @"Vl�@cY���#Z�b�tyE3�8S����@,"Vl�@�%|���@��bS�D�q ~ q ~       q ~ sq ~ @"Vl�@cY���#Z�b�N�k�d�7��%��@,"Vl�@�A]��I@���`�L'q ~ q ~       q ~ sq ~ @��D(\�@SY���#[�bE@�G���@�C� ^@#��D(\�@������@�[�ܤ9�q ~ q ~       q ~ sq ~ @��D(\�@SY���#[�bGͱҞ+�@����k@#��D(\�@�tY[��@�`���q ~ q ~       q ~ xpt player1q ~ pq ~ sq ~              �����  u                sq ~ @      @S��Y�C;                @$      @��     @x     sq ~     �  �pppq ~       q ~ sq ~     w   q ~ Zxpt player2q ~ [pq ~ x